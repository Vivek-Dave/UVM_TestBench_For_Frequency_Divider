`include "assertion_ip.sv"
`include "binding_module.sv"
`include "interface.sv"
`include "tb_pkg.sv"
module top;
  import uvm_pkg::*;
  import tb_pkg::*;
  
  bit clk; // external signal declaration

  //----------------------------------------------------------------------------
  intf i_intf(clk);
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  freq_divider DUT(.in(i_intf.in),
                   .clk(i_intf.clk),
                   .rst(i_intf.rst),
                   .out(i_intf.out)
                  );
  //----------------------------------------------------------------------------               
  
  initial begin
    clk<=0;
  end

  always #50 clk=~clk;
  
  //----------------------------------------------------------------------------
  initial begin
    $dumpfile("dumpfile.vcd");
    $dumpvars;
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    uvm_config_db#(virtual intf)::set(uvm_root::get(),"","vif",i_intf);
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    run_test("freq_div_test");
  end
  //----------------------------------------------------------------------------
endmodule

